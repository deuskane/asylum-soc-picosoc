-------------------------------------------------------------------------------
-- Title      : PicoSoC
-- Project    : 
-------------------------------------------------------------------------------
-- File       : PicoSoC.vhd
-- Author     : Mathieu Rosiere
-- Company    : 
-- Created    : 2017-03-30
-- Last update: 2025-12-03
-- Platform   : 
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: 
-------------------------------------------------------------------------------
-- Copyright (c) 2017 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author   Description
-- 2017-03-30  1.0      mrosiere Created
-- 2024-12-31  1.1      mrosiere Fix parameter to GPIO
-- 2025-01-12  2.0      mrosiere Add Safety feature
-- 2025-01-15  2.1      mrosiere Update diff detection
-- 2025-01-21  2.2      mrosiere Add UART
-- 2025-04-02  2.3      mrosiere Use ICN
-- 2025-07-15  3.0      mrosiere Add FIFO depth for UART and SPI
-- 2025-11-02  3.1      mrosiere Add Timer
-- 2025-11-27  3.2      mrosiere Add CRC
-- 2025-11-29  3.3      mrosiere Use CRC Generic
-------------------------------------------------------------------------------

library ieee;
use     ieee.std_logic_1164.all;
use     ieee.numeric_std.all;
library asylum;

-- CSR Package
use     asylum.GPIO_csr_pkg.all;
use     asylum.UART_csr_pkg.all;
use     asylum.SPI_csr_pkg.all;
use     asylum.GIC_csr_pkg.all;
use     asylum.timer_csr_pkg.all;
use     asylum.crc_csr_pkg.all;
-- Type Package
use     asylum.sbi_pkg.all;
-- Modules Packages
use     asylum.PicoSoC_pkg.all;
use     asylum.OpenBlaze8_pkg.all;
use     asylum.gpio_pkg.all;
use     asylum.uart_pkg.all;
use     asylum.spi_pkg.all;
use     asylum.gic_pkg.all;
use     asylum.timer_pkg.all;
use     asylum.crc_pkg.all;
use     asylum.icn_pkg.all;

entity PicoSoC_user is
  generic
    (CLOCK_FREQ            : integer  := 50000000
    ;BAUD_RATE             : integer  := 115200
    ;UART_DEPTH_TX         : natural  := 0
    ;UART_DEPTH_RX         : natural  := 0
    ;SPI_DEPTH_CMD         : natural  := 0
    ;SPI_DEPTH_TX          : natural  := 0
    ;SPI_DEPTH_RX          : natural  := 0
    ;NB_SWITCH             : positive := 8
    ;NB_LED0               : positive := 8
    ;NB_LED1               : positive := 8
    ;SAFETY                : string   := "lock-step" -- "none" / "lock-step" / "tmr"
    ;FAULT_INJECTION       : boolean  := False
    
    ;ICN_ALGO_SEL          : string := "or"
    );
  port
    (clk_i                 : in  std_logic
    ;arst_b_i              : in  std_logic
                          
    ;switch_i              : in  std_logic_vector(NB_SWITCH-1 downto 0)
    ;led0_o                : out std_logic_vector(NB_LED0  -1 downto 0)
    ;led1_o                : out std_logic_vector(NB_LED1  -1 downto 0)

     -- UART Interface
    ;uart_tx_o             : out std_logic
    ;uart_rx_i             : in  std_logic
    ;uart_cts_b_i          : in  std_logic -- Clear   To Send (Active low)
    ;uart_rts_b_o          : out std_logic -- Request To Send (Active low)
                          
    -- SPI Interface
    ;spi_sclk_o            : out std_logic
    ;spi_cs_b_o            : out std_logic
    ;spi_mosi_o            : out std_logic
    ;spi_miso_i            : in  std_logic
                          
    ;it_i                  : in  std_logic
    ;inject_error_i        : in  std_logic_vector(        3-1 downto 0)
    ;diff_o                : out std_logic_vector(        3-1 downto 0) -- bit 0 : cpu0 vs cpu1
                                                                        -- bit 1 : cpu1 vs cpu2
                                                                        -- bit 2 : cpu2 vs cpu0
                                 
    ;debug_o               : out PicoSoC_user_debug_t
    );
end PicoSoC_user;

architecture rtl of PicoSoC_user is

  -- Constant declaration
  constant CST0                       : std_logic_vector (8-1 downto 0) := (others => '0');
  constant CST1                       : std_logic_vector (8-1 downto 0) := (others => '1');

  -- Module parameters
  constant CPU1_ENABLE                : boolean := ((SAFETY = "lock-step") or
                                                    (SAFETY = "tmr"));
  constant CPU2_ENABLE                : boolean := ((SAFETY = "tmr"));

  -- ICN Configuration
  constant TARGET_ADDR_ENCODING       : string := PICOSOC_USER_ADDR_ENCODING;
  
  constant TARGET_SWITCH              : integer  := 0;
  constant TARGET_LED0                : integer  := 1;
  constant TARGET_LED1                : integer  := 2;
  constant TARGET_UART                : integer  := 3;
  constant TARGET_SPI                 : integer  := 4;
  constant TARGET_GIC                 : integer  := 5;
  constant TARGET_TIMER               : integer  := 6;
  constant TARGET_CRC                 : integer  := 7;
  
  constant NB_TARGET                  : positive := 8;
  
  constant TARGET_ID                  : sbi_addrs_t   (NB_TARGET-1 downto 0) :=
    ( TARGET_SWITCH                   => PICOSOC_USER_SWITCH_BA
     ,TARGET_LED0                     => PICOSOC_USER_LED0_BA  
     ,TARGET_LED1                     => PICOSOC_USER_LED1_BA  
     ,TARGET_UART                     => PICOSOC_USER_UART_BA  
     ,TARGET_SPI                      => PICOSOC_USER_SPI_BA   
     ,TARGET_GIC                      => PICOSOC_USER_GIC_BA   
     ,TARGET_TIMER                    => PICOSOC_USER_TIMER_BA 
     ,TARGET_CRC                      => PICOSOC_USER_CRC_BA   
      );

  constant TARGET_ADDR_WIDTH          : naturals_t    (NB_TARGET-1 downto 0) :=
    ( TARGET_SWITCH                   => GPIO_ADDR_WIDTH
     ,TARGET_LED0                     => GPIO_ADDR_WIDTH
     ,TARGET_LED1                     => GPIO_ADDR_WIDTH
     ,TARGET_UART                     => UART_ADDR_WIDTH
     ,TARGET_SPI                      => SPI_ADDR_WIDTH
     ,TARGET_GIC                      => GIC_ADDR_WIDTH
     ,TARGET_TIMER                    => TIMER_ADDR_WIDTH
     ,TARGET_CRC                      => CRC_ADDR_WIDTH
      );
  
  -- Signals ICN
  signal   icn_sbi_inis               : sbi_inis_t(NB_TARGET-1 downto 0)(addr (SBI_ADDR_WIDTH-1 downto 0),
                                                                         wdata(SBI_DATA_WIDTH-1 downto 0));
  signal   icn_sbi_tgts               : sbi_tgts_t(NB_TARGET-1 downto 0)(rdata(SBI_DATA_WIDTH-1 downto 0));

  -- Signals Clock/Reset
  signal   clk                        : std_logic;
  signal   arst_b                     : std_logic;

  -- Signals CPUs
  signal   cpu0_ics                   : std_logic;
  signal   cpu0_iaddr                 : std_logic_vector(10-1 downto 0);
  signal   cpu0_idata                 : std_logic_vector(18-1 downto 0);
  signal   cpu0_sbi_ini               : sbi_ini_t(addr (SBI_ADDR_WIDTH-1 downto 0),
                                                  wdata(SBI_DATA_WIDTH-1 downto 0));
  signal   cpu0_it_ack                : std_logic;
  
  signal   cpu1_ics                   : std_logic;
  signal   cpu1_iaddr                 : std_logic_vector(10-1 downto 0);
  signal   cpu1_idata                 : std_logic_vector(18-1 downto 0);
  signal   cpu1_sbi_ini               : sbi_ini_t(addr (SBI_ADDR_WIDTH-1 downto 0),
                                                  wdata(SBI_DATA_WIDTH-1 downto 0));
  signal   cpu1_it_ack                : std_logic;
  
  signal   cpu2_ics                   : std_logic;
  signal   cpu2_iaddr                 : std_logic_vector(10-1 downto 0);
  signal   cpu2_idata                 : std_logic_vector(18-1 downto 0);
  signal   cpu2_sbi_ini               : sbi_ini_t(addr (SBI_ADDR_WIDTH-1 downto 0),
                                                  wdata(SBI_DATA_WIDTH-1 downto 0));
  signal   cpu2_it_ack                : std_logic;

  -- Signals CPU (post lockstep / TMR)
  signal   cpu_ics                    : std_logic;
  signal   cpu_iaddr                  : std_logic_vector(10-1 downto 0);
  signal   cpu_idata                  : std_logic_vector(18-1 downto 0);

  signal   cpu_sbi_ini                : sbi_ini_t(addr (SBI_ADDR_WIDTH-1 downto 0),
                                                  wdata(SBI_DATA_WIDTH-1 downto 0));
  signal   cpu_sbi_tgt                : sbi_tgt_t(rdata(SBI_DATA_WIDTH-1 downto 0));
  signal   cpu_it_val                 : std_logic;
  signal   cpu_it_ack                 : std_logic;

  -- UART
  signal   uart_it                    : std_logic;
  
  -- Interruption Vector

  constant GIC_IT_USER                : natural  := 0;
  constant GIC_UART                   : natural  := 1;
  constant GIC_TIMER                  : natural  := 2;

  constant GIC_WIDTH                  : positive := 3;

  signal   gic_it_vector              : std_logic_vector(GIC_WIDTH-1 downto 0);

  -- Timer
  signal   timer_disable              : std_logic;
  signal   timer_clear                : std_logic;
  signal   timer_it                   : std_logic;
  
  -- Signals Safety
  signal   diff                       : std_logic_vector(3-1 downto 0); -- bit 0 : cpu0 vs cpu1
                                                                        -- bit 1 : cpu1 vs cpu2
                                                                        -- bit 2 : cpu2 vs cpu0
  signal   diff_r                     : std_logic_vector(3-1 downto 0); -- bit 0 : cpu0 vs cpu1
                                                                        -- bit 1 : cpu1 vs cpu2
                                                                        -- bit 2 : cpu2 vs cpu0

begin  -- architecture rtl

  -----------------------------------------------------------------------------
  -- Clock & Reset
  -----------------------------------------------------------------------------
  clk    <= clk_i;
  arst_b <= arst_b_i;
  
  -----------------------------------------------------------------------------
  -- CPU 0
  -----------------------------------------------------------------------------
  ins_sbi_OpenBlaze8_0 : sbi_OpenBlaze8
    generic map
    (RAM_DEPTH            => 256,
     REGFILE_SYNC_READ    => true
     )
    port map
    (clk_i                => clk         
    ,cke_i                => '1'         
    ,arstn_i              => arst_b      
    ,ics_o                => cpu0_ics    
    ,iaddr_o              => cpu0_iaddr  
    ,idata_i              => cpu0_idata  
    ,sbi_ini_o            => cpu0_sbi_ini
    ,sbi_tgt_i            => cpu_sbi_tgt 
    ,interrupt_i          => cpu_it_val  
    ,interrupt_ack_o      => cpu0_it_ack
    );

  -----------------------------------------------------------------------------
  -- CPU ROM
  -----------------------------------------------------------------------------
  ins_sbi_OpenBlaze8_ROM : entity asylum.ROM_user(rom)
    port map
    (clk_i                => clk      
    ,cke_i                => cpu_ics  
    ,address_i            => cpu_iaddr
    ,instruction_o        => cpu_idata
    );

  -----------------------------------------------------------------------------
  -- CPU Signals
  --  * ROM interface
  --  * ICN interface
  --  * IT  interface
  --
  -- If safety none or lock-step : take cpu 0
  -- else if tmr : vote all cpu output
  -----------------------------------------------------------------------------
  gen_cpu_vote: if SAFETY = "tmr"
  generate
    cpu_ics        <= ((cpu0_ics     and cpu1_ics    ) or
                       (cpu1_ics     and cpu2_ics    ) or
                       (cpu2_ics     and cpu0_ics    ));
    cpu_iaddr      <= ((cpu0_iaddr   and cpu1_iaddr  ) or
                       (cpu1_iaddr   and cpu2_iaddr  ) or
                       (cpu2_iaddr   and cpu0_iaddr  ));
    cpu_sbi_ini    <= ((cpu0_sbi_ini and cpu1_sbi_ini) or
                       (cpu1_sbi_ini and cpu2_sbi_ini) or
                       (cpu2_sbi_ini and cpu0_sbi_ini));
    cpu_it_ack     <= ((cpu0_it_ack  and cpu1_it_ack ) or
                       (cpu1_it_ack  and cpu2_it_ack ) or
                       (cpu2_it_ack  and cpu0_it_ack ));
  end generate;

  gen_cpu_vote_b: if SAFETY /= "tmr"
  generate
    cpu_ics        <= cpu0_ics     ;
    cpu_iaddr      <= cpu0_iaddr   ;
    cpu_sbi_ini    <= cpu0_sbi_ini ;
    cpu_it_ack     <= cpu0_it_ack  ;
  end generate;
  
  -----------------------------------------------------------------------------
  -- Interconnect
  -- From 1 Initiator to N Target
  -----------------------------------------------------------------------------
  ins_sbi_icn : sbi_icn
    generic map
    (NB_TARGET            => NB_TARGET
    ,TARGET_ID            => TARGET_ID
    ,TARGET_ADDR_WIDTH    => TARGET_ADDR_WIDTH
    ,TARGET_ADDR_ENCODING => TARGET_ADDR_ENCODING
    ,ALGO_SEL             => ICN_ALGO_SEL
      )
    port map
    (clk_i                => clk      
    ,cke_i                => '1'         
    ,arst_b_i             => arst_b      
    ,sbi_ini_i            => cpu_sbi_ini 
    ,sbi_tgt_o            => cpu_sbi_tgt 
    ,sbi_inis_o           => icn_sbi_inis
    ,sbi_tgts_i           => icn_sbi_tgts
    );

  -----------------------------------------------------------------------------
  -- GPIO 0 - Switch
  -----------------------------------------------------------------------------
  ins_sbi_switch : sbi_GPIO
    generic map
    (NB_IO                => NB_SWITCH
    ,DATA_OE_INIT         => CST0(8-1 downto 0)
    ,IT_ENABLE            => false
    )
    port map
    (clk_i                => clk           
    ,cke_i                => '1'           
    ,arstn_i              => arst_b         
    ,sbi_ini_i            => icn_sbi_inis(TARGET_SWITCH)   
    ,sbi_tgt_o            => icn_sbi_tgts(TARGET_SWITCH)   
    ,data_i               => switch_i      
    ,data_o               => open          
    ,data_oe_o            => open          
    ,interrupt_o          => open          
    ,interrupt_ack_i      => '0'
    );

  -----------------------------------------------------------------------------
  -- GPIO 1 - LED
  -----------------------------------------------------------------------------
  ins_sbi_led0 : sbi_GPIO
    generic map
    (NB_IO                => NB_LED0
    ,DATA_OE_INIT         => CST1(8-1 downto 0)
    ,IT_ENABLE            => false
    )
    port map
    (clk_i                => clk         
    ,cke_i                => '1'         
    ,arstn_i              => arst_b       
    ,sbi_ini_i            => icn_sbi_inis(TARGET_LED0) 
    ,sbi_tgt_o            => icn_sbi_tgts(TARGET_LED0) 
    ,data_i               => X"00"       
    ,data_o               => led0_o      
    ,data_oe_o            => open        
    ,interrupt_o          => open        
    ,interrupt_ack_i      => '0'
    );

  -----------------------------------------------------------------------------
  -- GPIO 2 - LED
  -----------------------------------------------------------------------------
  ins_sbi_led1 : sbi_GPIO
    generic map
    (NB_IO                => NB_LED1
    ,DATA_OE_INIT         => CST1(8-1 downto 0)
    ,IT_ENABLE            => false
    )
    port map
    (clk_i                => clk         
    ,cke_i                => '1'         
    ,arstn_i              => arst_b       
    ,sbi_ini_i            => icn_sbi_inis(TARGET_LED1) 
    ,sbi_tgt_o            => icn_sbi_tgts(TARGET_LED1) 
    ,data_i               => X"00"       
    ,data_o               => led1_o      
    ,data_oe_o            => open        
    ,interrupt_o          => open        
    ,interrupt_ack_i      => '0'
    );

  -----------------------------------------------------------------------------
  -- UART
  -----------------------------------------------------------------------------
  ins_sbi_uart : sbi_uart
    generic map
    (BAUD_RATE            => BAUD_RATE     
    ,CLOCK_FREQ           => CLOCK_FREQ
    ,DEPTH_TX             => UART_DEPTH_TX 
    ,DEPTH_RX             => UART_DEPTH_RX 
     )
    port map
    (clk_i                => clk           
    ,arst_b_i             => arst_b        
    ,sbi_ini_i            => icn_sbi_inis(TARGET_UART)   
    ,sbi_tgt_o            => icn_sbi_tgts(TARGET_UART)   
    ,uart_tx_o            => uart_tx_o     
    ,uart_rx_i            => uart_rx_i
    ,uart_cts_b_i         => uart_cts_b_i
    ,uart_rts_b_o         => uart_rts_b_o
    ,it_o                 => uart_it
    ,debug_o              => debug_o.uart
     );

  -----------------------------------------------------------------------------
  -- SPI
  -----------------------------------------------------------------------------
  ins_sbi_spi : sbi_spi
    generic map
    (USER_DEFINE_PRESCALER=> true
    ,PRESCALER_RATIO      => x"00"
    ,DEPTH_CMD            => SPI_DEPTH_CMD
    ,DEPTH_TX             => SPI_DEPTH_TX 
    ,DEPTH_RX             => SPI_DEPTH_RX 
     )
    port map
    (clk_i                => clk           
    ,arst_b_i             => arst_b        
    ,sbi_ini_i            => icn_sbi_inis(TARGET_SPI)   
    ,sbi_tgt_o            => icn_sbi_tgts(TARGET_SPI)   
    ,sclk_o               => spi_sclk_o   
    ,sclk_oe_o            => open
    ,cs_b_o               => spi_cs_b_o   
    ,cs_b_oe_o            => open
    ,mosi_o               => spi_mosi_o   
    ,mosi_oe_o            => open
    ,miso_i               => spi_miso_i   
     );

  -----------------------------------------------------------------------------
  -- GIC - Interruption Vector
  -----------------------------------------------------------------------------
  gic_it_vector(GIC_IT_USER) <= it_i   ;
  gic_it_vector(GIC_UART   ) <= uart_it;
  gic_it_vector(GIC_TIMER  ) <= timer_it;

  ins_sbi_gic : sbi_GIC
    port map
    (clk_i                => clk         
    ,arst_b_i             => arst_b      
    ,sbi_ini_i            => icn_sbi_inis(TARGET_GIC)
    ,sbi_tgt_o            => icn_sbi_tgts(TARGET_GIC)
    ,its_i                => gic_it_vector
    ,itm_o                => cpu_it_val
    );

  -----------------------------------------------------------------------------
  -- Timer
  -----------------------------------------------------------------------------
  timer_disable <= '0';
  timer_clear   <= '0';

  ins_sbi_timer : sbi_timer
    port map
    (clk_i                => clk         
    ,arst_b_i             => arst_b      
    ,sbi_ini_i            => icn_sbi_inis(TARGET_TIMER)
    ,sbi_tgt_o            => icn_sbi_tgts(TARGET_TIMER)
    ,timer_disable_i      => timer_disable
    ,timer_clear_i        => timer_clear
    ,it_o                 => timer_it
    );
  
  -----------------------------------------------------------------------------
  -- CRC
  -----------------------------------------------------------------------------
  ins_sbi_crc : sbi_crc
    generic map
    (WIDTH_CRC        => 16      ,
     WIDTH_DATA       => 8       ,
     POLYNOM          => X"A001" ,
     SHIFT_LEFT       => false   ,
     LSB_FIRST        => true    ,
     POLYNOM_REVERSE  => false   ,
     REFLECT_IN       => false   ,
     REFLECT_OUT      => false   ,
     XOR_OUT          => (others => '0')
      )
    port map
    (clk_i                => clk         
    ,arst_b_i             => arst_b      
    ,sbi_ini_i            => icn_sbi_inis(TARGET_CRC)
    ,sbi_tgt_o            => icn_sbi_tgts(TARGET_CRC)
    );

  -----------------------------------------------------------------------------
  -- CPU 1
  -- diff cpu0 vs cpu1
  -----------------------------------------------------------------------------
  gen_cpu1_enable: if CPU1_ENABLE = true
  generate
    -- Lock Step
    ins_sbi_OpenBlaze8_1 : sbi_OpenBlaze8
      generic map
      (RAM_DEPTH            => 256,
       REGFILE_SYNC_READ    => true
       )
      port map
      (clk_i                => clk           
      ,cke_i                => '1'     
      ,arstn_i              => arst_b   
      ,ics_o                => cpu1_ics    
      ,iaddr_o              => cpu1_iaddr  
      ,idata_i              => cpu1_idata  
      ,sbi_ini_o            => cpu1_sbi_ini
      ,sbi_tgt_i            => cpu_sbi_tgt 
      ,interrupt_i          => cpu_it_val  
      ,interrupt_ack_o      => cpu1_it_ack
       );

    diff(0) <= '1' when (   (cpu0_ics           /= cpu1_ics          )
                         or (cpu0_iaddr         /= cpu1_iaddr        )
                         or (cpu0_it_ack        /= cpu1_it_ack       )
                       --or (cpu0_sbi_ini       /= cpu1_sbi_ini      )
                            ) else
               '0';
    
    p_diff_r: process (clk, arst_b) is
    begin  -- process p_diff_r
      if arst_b = '0' then                 -- asynchronous reset (active low)
        diff_r(0) <= '0';
      elsif clk'event and clk = '1' then  -- rising clock edge
        -- Trap 1
        diff_r(0) <= diff_r(0) or diff(0);
      end if;
    end process p_diff_r;

    diff_o(0) <= diff_r(0);
  end generate gen_cpu1_enable;
  
  gen_cpu1_disable: if CPU1_ENABLE = false
  generate
    diff_o(0) <= '0';
  end generate gen_cpu1_disable;

  -----------------------------------------------------------------------------
  -- CPU 2
  -- diff cpu1 vs cpu2
  -- diff cpu2 vs cpu0
  -----------------------------------------------------------------------------
  gen_cpu2_enable: if CPU2_ENABLE = true
  generate
    -- TMR
    ins_sbi_OpenBlaze8_2 : sbi_OpenBlaze8
      generic map
      (RAM_DEPTH            => 256,
       REGFILE_SYNC_READ    => true
       )
      port map
      (clk_i                => clk           
      ,cke_i                => '1'     
      ,arstn_i              => arst_b   
      ,ics_o                => cpu2_ics    
      ,iaddr_o              => cpu2_iaddr  
      ,idata_i              => cpu2_idata  
      ,sbi_ini_o            => cpu2_sbi_ini
      ,sbi_tgt_i            => cpu_sbi_tgt 
      ,interrupt_i          => cpu_it_val  
      ,interrupt_ack_o      => cpu2_it_ack
       );

    diff(1) <= '1' when (   (cpu1_ics           /= cpu2_ics          )
                         or (cpu1_iaddr         /= cpu2_iaddr        )
                         or (cpu1_it_ack        /= cpu2_it_ack       )
                       --or (cpu1_sbi_ini       /= cpu2_sbi_ini      )
                         ) else
               '0';
    diff(2) <= '1' when (   (cpu2_ics           /= cpu0_ics          )
                         or (cpu2_iaddr         /= cpu0_iaddr        )
                         or (cpu2_it_ack        /= cpu0_it_ack       )
                       --or (cpu2_sbi_ini       /= cpu0_sbi_ini      )
                         ) else
               '0';
    
    p_diff_r: process (clk, arst_b) is
    begin  -- process p_diff_r
      if arst_b = '0' then                 -- asynchronous reset (active low)
        diff_r(2 downto 1) <= "00";
      elsif clk'event and clk = '1' then  -- rising clock edge

        -- Trap 1
        diff_r(2 downto 1) <= diff_r(2 downto 1) or diff(2 downto 1);
      end if;
    end process p_diff_r;

    diff_o(2 downto 1) <= diff_r(2 downto 1);
  end generate gen_cpu2_enable;
  
  gen_cpu2_disable: if CPU2_ENABLE = false
  generate
    diff_o(1) <= '0';
    diff_o(2) <= '0';
  end generate gen_cpu2_disable;

  -----------------------------------------------------------------------------
  -- Fault Injection
  -----------------------------------------------------------------------------
  gen_inject_error:   if FAULT_INJECTION = true
  generate
    cpu0_idata(17)          <= cpu_idata(17) xor inject_error_i(0);
    cpu0_idata(16 downto 0) <= cpu_idata(16 downto 0);

    cpu1_idata(17)          <= cpu_idata(17) xor inject_error_i(1);
    cpu1_idata(16 downto 0) <= cpu_idata(16 downto 0);

    cpu2_idata(17)          <= cpu_idata(17) xor inject_error_i(2);
    cpu2_idata(16 downto 0) <= cpu_idata(16 downto 0);
        
  end generate gen_inject_error;

  gen_inject_error_n: if FAULT_INJECTION = false
  generate
    cpu0_idata              <= cpu_idata;
    cpu1_idata              <= cpu_idata;        
    cpu2_idata              <= cpu_idata;        
  end generate gen_inject_error_n;

  -----------------------------------------------------------------------------
  -- Debug
  -----------------------------------------------------------------------------
  debug_o.arst_b      <= arst_b                           ;
  debug_o.cpu_iaddr   <= cpu_iaddr                        ;
  debug_o.cpu_idata   <= cpu_idata                        ;
  debug_o.cpu_dcs     <= cpu_sbi_ini.cs                   ;
  debug_o.cpu_dre     <= cpu_sbi_ini.re                   ;
  debug_o.cpu_dwe     <= cpu_sbi_ini.we                   ;
  debug_o.cpu_daddr   <= cpu_sbi_ini.addr                 ;
  debug_o.cpu_dready  <= cpu_sbi_tgt.ready                ;
  debug_o.switch_cs   <= icn_sbi_inis(TARGET_SWITCH).cs   ;
  debug_o.switch_ready<= icn_sbi_tgts(TARGET_SWITCH).ready;
  debug_o.led0_cs     <= icn_sbi_inis(TARGET_LED0  ).cs   ;
  debug_o.led0_ready  <= icn_sbi_tgts(TARGET_LED0  ).ready;
  debug_o.led1_cs     <= icn_sbi_inis(TARGET_LED1  ).cs   ;
  debug_o.led1_ready  <= icn_sbi_tgts(TARGET_LED1  ).ready;
  debug_o.uart_cs     <= icn_sbi_inis(TARGET_UART  ).cs   ;
  debug_o.uart_ready  <= icn_sbi_tgts(TARGET_UART  ).ready;
  debug_o.spi_cs      <= icn_sbi_inis(TARGET_SPI   ).cs   ;
  debug_o.spi_ready   <= icn_sbi_tgts(TARGET_SPI   ).ready;
    
end architecture rtl;
    
